module a_and_b (
    input       a,
    input       b,
    output      c
);

and (c,a,b);
    
endmodule